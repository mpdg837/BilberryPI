	module KERNAL(
       input clk,
       input[11:0] addr,
       output reg[31:0] out
);

wire[31:0] out1;
wire[31:0] out2;
wire[31:0] out3;

ROM1 r1(.clk(clk),
     .addr(addr),
     .out(out1)
);

ROM2 r2(.clk(clk),
     .addr(addr+1024),
     .out(out2)
);

reg[1:0] bufstat;

always@(posedge clk)begin
	bufstat <= addr[10:9];
end

always@(*)begin
	case(bufstat)
		0: out= out1;
		1: out= out1;
		2: out= out2;
		3: out= out2;
	endcase
end

endmodule

module ROM1(
       input clk,
       input[11:0] addr,
       output reg[31:0] out
);

always@(posedge clk)
case(addr[9:0])
11'd0: out <= 32'b00000001111100000000000000000001;
11'd1: out <= 32'b00000000010100000000000010011110;
11'd2: out <= 32'b00000000010100000000000001001011;
11'd3: out <= 32'b00000000010100000000001000100110;
11'd4: out <= 32'b00000000010100000000000000111100;
11'd5: out <= 32'b00000000010100000000000101000110;
11'd6: out <= 32'b00000000010100000000000101010001;
11'd7: out <= 32'b00000000010100000000001000111100;
11'd8: out <= 32'b00000000010100000000000011011101;
11'd9: out <= 32'b00000000000100000000000000000000;
11'd10: out <= 32'b00000000000101000000000000000000;
11'd11: out <= 32'b00000000000110000000000000000000;
11'd12: out <= 32'b00000000000111000000000000000000;
11'd13: out <= 32'b00000001111100000000000000000000;
11'd14: out <= 32'b00000001101100000000000000000000;
11'd15: out <= 32'b00000000011000000000000000000000;
11'd16: out <= 32'b00000001101100000000000000000000;
11'd17: out <= 32'b00000000011001000000000000000000;
11'd18: out <= 32'b00000001101100000000000000000000;
11'd19: out <= 32'b00000000011010000000000000000000;
11'd20: out <= 32'b00000001101100000000000000000000;
11'd21: out <= 32'b00000000011011000000000000000000;
11'd22: out <= 32'b00000001111100000000000000000000;
11'd23: out <= 32'b00000001111000000000000000001110;
11'd24: out <= 32'b00000001111000000000000000001001;
11'd25: out <= 32'b00000001111100000000000000000000;
11'd26: out <= 32'b00000000011100000001111111110100;
11'd27: out <= 32'b00000000011000000000000000000000;
11'd28: out <= 32'b00000000011100000001111111110101;
11'd29: out <= 32'b00000000011001000000000000000000;
11'd30: out <= 32'b00000000011100000001111111110110;
11'd31: out <= 32'b00000000011010000000000000000000;
11'd32: out <= 32'b00000000011100000001111111110111;
11'd33: out <= 32'b00000000011011000000000000000000;
11'd34: out <= 32'b00000001111000000000000000001001;
11'd35: out <= 32'b00000001111100000000000000000000;
11'd36: out <= 32'b00000001101000000000000000000000;
11'd37: out <= 32'b00000001100011000000000000000000;
11'd38: out <= 32'b00000001101000000000000000000000;
11'd39: out <= 32'b00000001100010000000000000000000;
11'd40: out <= 32'b00000001101000000000000000000000;
11'd41: out <= 32'b00000001100001000000000000000000;
11'd42: out <= 32'b00000001101000000000000000000000;
11'd43: out <= 32'b00000001100000000000000000000000;
11'd44: out <= 32'b00000001111100000000000000000000;
11'd45: out <= 32'b00000000011100000001111111110100;
11'd46: out <= 32'b00000001100000000000000000000000;
11'd47: out <= 32'b00000000011100000001111111110101;
11'd48: out <= 32'b00000001100001000000000000000000;
11'd49: out <= 32'b00000000011100000001111111110110;
11'd50: out <= 32'b00000001100010000000000000000000;
11'd51: out <= 32'b00000000011100000001111111110111;
11'd52: out <= 32'b00000001100011000000000000000000;
11'd53: out <= 32'b00000001111100000000000000000000;
11'd54: out <= 32'b00000001111000000000000000001110;
11'd55: out <= 32'b00000000111000000100000000000000;
11'd56: out <= 32'b00000000001101000000000000000000;
11'd57: out <= 32'b00000000001100000000000000000001;
11'd58: out <= 32'b00000001111000000000000000100100;
11'd59: out <= 32'b00000001111100000000000000000000;
11'd60: out <= 32'b00000001111000000000000000011010;
11'd61: out <= 32'b00000000000011000000000000000001;
11'd62: out <= 32'b00000000001000000000000000000000;
11'd63: out <= 32'b00000000110100001000000000000000;
11'd64: out <= 32'b00000001011100001000000000000000;
11'd65: out <= 32'b00000001001000000000000001000110;
11'd66: out <= 32'b00000000001000000000000000000000;
11'd67: out <= 32'b00000000011100000010000100011111;
11'd68: out <= 32'b00000000011000000000000000000000;
11'd69: out <= 32'b00000000010100000000000001001001;
11'd70: out <= 32'b00000000001000000000000000000000;
11'd71: out <= 32'b00000000011100000010000100011110;
11'd72: out <= 32'b00000000011000000000000000000000;
11'd73: out <= 32'b00000001111000000000000000101101;
11'd74: out <= 32'b00000001111100000000000000000000;
11'd75: out <= 32'b00000001111000000000000000011010;
11'd76: out <= 32'b00000000011100000010000100010001;
11'd77: out <= 32'b00000001100000000000000000000000;
11'd78: out <= 32'b00000001011100001111111111111111;
11'd79: out <= 32'b00000001001000000000000001010110;
11'd80: out <= 32'b00000000000011000000000000000010;
11'd81: out <= 32'b00000000001000000000000000000000;
11'd82: out <= 32'b00000000110100000000000000001111;
11'd83: out <= 32'b00000000011100000001111111100000;
11'd84: out <= 32'b00000000011000000000000000000000;
11'd85: out <= 32'b00000001111000000000000100001110;
11'd86: out <= 32'b00000001111000000000000000101101;
11'd87: out <= 32'b00000001111100000000000000000000;
11'd88: out <= 32'b00000000010100000000000001011000;
11'd89: out <= 32'b00000000100100000000000000000000;
11'd90: out <= 32'b00000000011011000000000000000000;
11'd91: out <= 32'b00000000011100000001000000000000;
11'd92: out <= 32'b00000000100100000000000000000000;
11'd93: out <= 32'b00000001100001000000000000000000;
11'd94: out <= 32'b00000001011101110000000000000000;
11'd95: out <= 32'b00000001001000000000000001100001;
11'd96: out <= 32'b00000000010100000000000001011000;
11'd97: out <= 32'b00000001111100000000000000000000;
11'd98: out <= 32'b00000000000100000001000000000000;
11'd99: out <= 32'b00000000000111000000000000000000;
11'd100: out <= 32'b00000001111000000000000001011001;
11'd101: out <= 32'b00000000010000000000000000000000;
11'd102: out <= 32'b00000001011100000011000000000000;
11'd103: out <= 32'b00000001001000000000000001101001;
11'd104: out <= 32'b00000000010100000000000001100011;
11'd105: out <= 32'b00000001111000000000000000001001;
11'd106: out <= 32'b00000001111100000000000000000000;
11'd107: out <= 32'b00000000000100000000000000001101;
11'd108: out <= 32'b00000000011100000010000100001010;
11'd109: out <= 32'b00000001100001000000000000000000;
11'd110: out <= 32'b00000001111000000000000100100000;
11'd111: out <= 32'b00000001111100000000000000000000;
11'd112: out <= 32'b00000001011100000000000000000000;
11'd113: out <= 32'b00000001010100000000000001110011;
11'd114: out <= 32'b00000000010100000000000001110101;
11'd115: out <= 32'b00000000101000000000000000000000;
11'd116: out <= 32'b00000000010000000000000000000000;
11'd117: out <= 32'b00000001111100000000000000000000;
11'd118: out <= 32'b00000001111000000000000000010111;
11'd119: out <= 32'b00000001111000000000001100111100;
11'd120: out <= 32'b00000000011100000001111111100001;
11'd121: out <= 32'b00000001100001000000000000000000;
11'd122: out <= 32'b00000001111000000000000100100000;
11'd123: out <= 32'b00000001111000000000000001101011;
11'd124: out <= 32'b00000001111000000000000000100100;
11'd125: out <= 32'b00000001111100000000000000000000;
11'd126: out <= 32'b00000001111000000000000000010111;
11'd127: out <= 32'b00000001111000000000001100111100;
11'd128: out <= 32'b00000000000101000000000000111110;
11'd129: out <= 32'b00000001111000000000000100100000;
11'd130: out <= 32'b00000001111000000000000001101011;
11'd131: out <= 32'b00000001111000000000000000100100;
11'd132: out <= 32'b00000001111100000000000000000000;
11'd133: out <= 32'b00000000011100000001111111000000;
11'd134: out <= 32'b00000000011000000000000000000000;
11'd135: out <= 32'b00000000011100000001111111000001;
11'd136: out <= 32'b00000000011001000000000000000000;
11'd137: out <= 32'b00000001111100000000000000000000;
11'd138: out <= 32'b00000001111000000000000001100010;
11'd139: out <= 32'b00000001111000000000000110010010;
11'd140: out <= 32'b00000001111000000000000110110001;
11'd141: out <= 32'b00000001111000000000000110101000;
11'd142: out <= 32'b00000001111000000000000111000001;
11'd143: out <= 32'b00000001111000000000000110101000;
11'd144: out <= 32'b00000001111000000000000111000001;
11'd145: out <= 32'b00000001111000000000000110101000;
11'd146: out <= 32'b00000001111000000000000111000001;
11'd147: out <= 32'b00000001111000000000000110101000;
11'd148: out <= 32'b00000001111000000000000111000001;
11'd149: out <= 32'b00000001111100000000000000000000;
11'd150: out <= 32'b00000001111000000000000010001010;
11'd151: out <= 32'b00000000000100000000000000000101;
11'd152: out <= 32'b00000000000101000000000000000000;
11'd153: out <= 32'b00000001111000000000000000110110;
11'd154: out <= 32'b00000000011100000010000100010000;
11'd155: out <= 32'b00000000011000000000100000000000;
11'd156: out <= 32'b00000001111000000000000101101101;
11'd157: out <= 32'b00000001111100000000000000000000;
11'd158: out <= 32'b00000001111000000000000010010110;
11'd159: out <= 32'b00000001111000000000001001010000;
11'd160: out <= 32'b00000001111000000000000010111100;
11'd161: out <= 32'b00000000000100000000000000000101;
11'd162: out <= 32'b00000000000101000000000000000010;
11'd163: out <= 32'b00000001111000000000000000110110;
11'd164: out <= 32'b00000000000100000000100000000010;
11'd165: out <= 32'b00000000010100000000000000000000;
11'd166: out <= 32'b00000001111000000000000000001110;
11'd167: out <= 32'b00000000011100000010000100010011;
11'd168: out <= 32'b00000000011000000001000000000000;
11'd169: out <= 32'b00000000011100000010000100011000;
11'd170: out <= 32'b00000001100001000000000000000000;
11'd171: out <= 32'b00000001101101000000000000000000;
11'd172: out <= 32'b00000000011001000000000000000000;
11'd173: out <= 32'b00000000011100000010000100011011;
11'd174: out <= 32'b00000001100000000000000000000000;
11'd175: out <= 32'b00000000011100000010000100011000;
11'd176: out <= 32'b00000000011000000000000000000000;
11'd177: out <= 32'b00000001111000000000000011000111;
11'd178: out <= 32'b00000001111000000000100000000010;
11'd179: out <= 32'b00000001101001000000000000000000;
11'd180: out <= 32'b00000001100001000000000000000000;
11'd181: out <= 32'b00000000011100000010000100011000;
11'd182: out <= 32'b00000000011001000000000000000000;
11'd183: out <= 32'b00000000011100000010000100010011;
11'd184: out <= 32'b00000000011000000001000000000000;
11'd185: out <= 32'b00000001111000000000000011000111;
11'd186: out <= 32'b00000001111000000000000000100100;
11'd187: out <= 32'b00000001111100000000000000000000;
11'd188: out <= 32'b00000001111000000000000000010111;
11'd189: out <= 32'b00000000011100000010000100010011;
11'd190: out <= 32'b00000000011000000001000000000000;
11'd191: out <= 32'b00000000011100000010000100011000;
11'd192: out <= 32'b00000000000100000000000000000000;
11'd193: out <= 32'b00000000011000000000000000000000;
11'd194: out <= 32'b00000000011100000010000100011011;
11'd195: out <= 32'b00000000011000000000000000000000;
11'd196: out <= 32'b00000001111000000000000011000111;
11'd197: out <= 32'b00000001111000000000000000100100;
11'd198: out <= 32'b00000001111100000000000000000000;
11'd199: out <= 32'b00000001111000000000000000001110;
11'd200: out <= 32'b00000001111000000000001001010101;
11'd201: out <= 32'b00000000011100000010000100010011;
11'd202: out <= 32'b00000001100000000000000000000000;
11'd203: out <= 32'b00000001011100000001001111111111;
11'd204: out <= 32'b00000001010000000000001010100011;
11'd205: out <= 32'b00000001001000000000001010100011;
11'd206: out <= 32'b00000000011100000010000100011000;
11'd207: out <= 32'b00000001100000000000000000000000;
11'd208: out <= 32'b00000000010000000000000000000000;
11'd209: out <= 32'b00000000011000000000000000000000;
11'd210: out <= 32'b00000000010100000000001010011000;
11'd211: out <= 32'b00000000011100000001000011111111;
11'd212: out <= 32'b00000001100000000000000000000000;
11'd213: out <= 32'b00000000011100000001111111100001;
11'd214: out <= 32'b00000000011000000000000000000000;
11'd215: out <= 32'b00000000011100000001011111111110;
11'd216: out <= 32'b00000000011000000000000001010000;
11'd217: out <= 32'b00000000011100000001011111111111;
11'd218: out <= 32'b00000000011000000001000000000000;
11'd219: out <= 32'b00000001111000000000000000100100;
11'd220: out <= 32'b00000001111100000000000000000000;
11'd221: out <= 32'b00000001111000000000000000011010;
11'd222: out <= 32'b00000000011100000010000100011100;
11'd223: out <= 32'b00000000011000001111111111111111;
11'd224: out <= 32'b00000000011100000010000100011101;
11'd225: out <= 32'b00000001100000000000000000000000;
11'd226: out <= 32'b00000001011100000111010100110000;
11'd227: out <= 32'b00000001001000000000000011100110;
11'd228: out <= 32'b00000000010000000000000000000000;
11'd229: out <= 32'b00000000011000000000000000000000;
11'd230: out <= 32'b00000001111000000000000000101101;
11'd231: out <= 32'b00000001111100000000000000000000;
11'd232: out <= 32'b00000001111000000000000000010111;
11'd233: out <= 32'b00000000011100000010000100011101;
11'd234: out <= 32'b00000000011000000000000000000000;
11'd235: out <= 32'b00000001111000000000000000100100;
11'd236: out <= 32'b00000001111100000000000000000000;
11'd237: out <= 32'b00000001111000000000000000001110;
11'd238: out <= 32'b00000000111000001111000000000000;
11'd239: out <= 32'b00000000001101000000000000000000;
11'd240: out <= 32'b00000000001100000000000000000001;
11'd241: out <= 32'b00000001111000000000000000100100;
11'd242: out <= 32'b00000001111100000000000000000000;
11'd243: out <= 32'b00000001111000000000000000010111;
11'd244: out <= 32'b00000000011100000010000000010000;
11'd245: out <= 32'b00000001100000000000000000000000;
11'd246: out <= 32'b00000001011100000000000000000000;
11'd247: out <= 32'b00000001001000000000000100000111;
11'd248: out <= 32'b00000000100100000000000000000000;
11'd249: out <= 32'b00000001100000000000000000000000;
11'd250: out <= 32'b00000001011100000000000011111111;
11'd251: out <= 32'b00000001001000000000000100000111;
11'd252: out <= 32'b00000000010100000000000011111101;
11'd253: out <= 32'b00000001100101000000000000000000;
11'd254: out <= 32'b00000000000100000000000000000001;
11'd255: out <= 32'b00000001111000000000000011101101;
11'd256: out <= 32'b00000000011100000010000000010000;
11'd257: out <= 32'b00000001100000000000000000000000;
11'd258: out <= 32'b00000000010000000000000000000000;
11'd259: out <= 32'b00000000011000000000000000000000;
11'd260: out <= 32'b00000000011100000010000000010001;
11'd261: out <= 32'b00000000011000001111111111111111;
11'd262: out <= 32'b00000000010100000000000100001100;
11'd263: out <= 32'b00000000011100000010000000010001;
11'd264: out <= 32'b00000000011000000000000000000000;
11'd265: out <= 32'b00000000000100000000000000000010;
11'd266: out <= 32'b00000000000101000000000000000000;
11'd267: out <= 32'b00000001111000000000000011101101;
11'd268: out <= 32'b00000001111000000000000000100100;
11'd269: out <= 32'b00000001111100000000000000000000;
11'd270: out <= 32'b00000000011100000001111111100000;
11'd271: out <= 32'b00000001100000000000000000000000;
11'd272: out <= 32'b00000000011100000010000100001000;
11'd273: out <= 32'b00000001100001000000000000000000;
11'd274: out <= 32'b00000001011100000000000000000001;
11'd275: out <= 32'b00000001001000000000000100010111;
11'd276: out <= 32'b00000001011100000000000000000010;
11'd277: out <= 32'b00000001001000000000000100011011;
11'd278: out <= 32'b00000000010100000000000100011111;
11'd279: out <= 32'b00000001011101010000000000000011;
11'd280: out <= 32'b00000001001000000000000100011111;
11'd281: out <= 32'b00000000010001000000000000000000;
11'd282: out <= 32'b00000000010100000000000100011110;
11'd283: out <= 32'b00000001011101010000000000000000;
11'd284: out <= 32'b00000001001000000000000100011110;
11'd285: out <= 32'b00000001011001000000000000000000;
11'd286: out <= 32'b00000000011001000000000000000000;
11'd287: out <= 32'b00000001111100000000000000000000;
11'd288: out <= 32'b00000001111000000000000000001110;
11'd289: out <= 32'b00000000111000001000000000000000;
11'd290: out <= 32'b00000000001101000000000000000000;
11'd291: out <= 32'b00000000001100000000000000000001;
11'd292: out <= 32'b00000001111000000000000000100100;
11'd293: out <= 32'b00000001111100000000000000000000;
11'd294: out <= 32'b00000001111000000000000000010111;
11'd295: out <= 32'b00000000011100000010000100000111;
11'd296: out <= 32'b00000001100011000000000000000000;
11'd297: out <= 32'b00000000000110000000000000000000;
11'd298: out <= 32'b00000000000100000000000000000011;
11'd299: out <= 32'b00000001100101100000000000000000;
11'd300: out <= 32'b00000001111000000000000100100000;
11'd301: out <= 32'b00000000000100000000000000000100;
11'd302: out <= 32'b00000000100111000000000000000000;
11'd303: out <= 32'b00000001100001000000000000000000;
11'd304: out <= 32'b00000001111000000000000100100000;
11'd305: out <= 32'b00000000010011000000000000000000;
11'd306: out <= 32'b00000000000100000000000000000101;
11'd307: out <= 32'b00000000100111000000000000000000;
11'd308: out <= 32'b00000001100001000000000000000000;
11'd309: out <= 32'b00000001111000000000000100100000;
11'd310: out <= 32'b00000000010011000000000000000000;
11'd311: out <= 32'b00000000010010000000000000000000;
11'd312: out <= 32'b00000001011110100000000000001000;
11'd313: out <= 32'b00000001001000000000000100111011;
11'd314: out <= 32'b00000000010100000000000100101010;
11'd315: out <= 32'b00000001111000000000000000100100;
11'd316: out <= 32'b00000001111100000000000000000000;
11'd317: out <= 32'b00000000000100000000000000000001;
11'd318: out <= 32'b00000000011100000010000100001101;
11'd319: out <= 32'b00000001100001000000000000000000;
11'd320: out <= 32'b00000001111000000000000100100000;
11'd321: out <= 32'b00000000000100000000000000000010;
11'd322: out <= 32'b00000000011100000010000100001110;
11'd323: out <= 32'b00000001100001000000000000000000;
11'd324: out <= 32'b00000001111000000000000100100000;
11'd325: out <= 32'b00000001111100000000000000000000;
11'd326: out <= 32'b00000001111100000000000000000010;
11'd327: out <= 32'b00000001111000000000000000011010;
11'd328: out <= 32'b00000000011100000010000100010001;
11'd329: out <= 32'b00000001100000000000000000000000;
11'd330: out <= 32'b00000001011100001111111111111111;
11'd331: out <= 32'b00000001001000000000000101001110;
11'd332: out <= 32'b00000000011100000001111111000010;
11'd333: out <= 32'b00000000011000001111111111111111;
11'd334: out <= 32'b00000001111100000000000000000001;
11'd335: out <= 32'b00000001111000000000000000101101;
11'd336: out <= 32'b00000001111100000000000000000000;
11'd337: out <= 32'b00000001111000000000000000011010;
11'd338: out <= 32'b00000000011100000010000000000010;
11'd339: out <= 32'b00000000011000001111111111111111;
11'd340: out <= 32'b00000001111000000000000000101101;
11'd341: out <= 32'b00000001111100000000000000000000;
11'd342: out <= 32'b00000001111000000000000000001110;
11'd343: out <= 32'b00000000000100000000000000010010;
11'd344: out <= 32'b00000001111000000000000100100000;
11'd345: out <= 32'b00000000000111000000000000000000;
11'd346: out <= 32'b00000000000100000000000000010011;
11'd347: out <= 32'b00000001100101110000000000000000;
11'd348: out <= 32'b00000001111000000000000100100000;
11'd349: out <= 32'b00000000100110000000000000000000;
11'd350: out <= 32'b00000001100001000000000000000000;
11'd351: out <= 32'b00000000000100000000000000010100;
11'd352: out <= 32'b00000001111000000000000100100000;
11'd353: out <= 32'b00000000010010000000000000000000;
11'd354: out <= 32'b00000000100110000000000000000000;
11'd355: out <= 32'b00000001100001000000000000000000;
11'd356: out <= 32'b00000000000100000000000000010101;
11'd357: out <= 32'b00000001111000000000000100100000;
11'd358: out <= 32'b00000000010010000000000000000000;
11'd359: out <= 32'b00000000010011000000000000000000;
11'd360: out <= 32'b00000001011111110000000000010000;
11'd361: out <= 32'b00000001001000000000000101101011;
11'd362: out <= 32'b00000000010100000000000101011010;
11'd363: out <= 32'b00000001111000000000000000100100;
11'd364: out <= 32'b00000001111100000000000000000000;
11'd365: out <= 32'b00000001111000000000000000001001;
11'd366: out <= 32'b00000000011100000010000100010000;
11'd367: out <= 32'b00000001100011000000000000000000;
11'd368: out <= 32'b00000000011100000010000100011001;
11'd369: out <= 32'b00000000000101000000000000000000;
11'd370: out <= 32'b00000000011001000000000000000000;
11'd371: out <= 32'b00000000011100000010000100011001;
11'd372: out <= 32'b00000001100001000000000000000000;
11'd373: out <= 32'b00000000000100000000000000000110;
11'd374: out <= 32'b00000001111000000000000100100000;
11'd375: out <= 32'b00000000000110000000000000000000;
11'd376: out <= 32'b00000000000100000000000000000111;
11'd377: out <= 32'b00000001100101100000000000000000;
11'd378: out <= 32'b00000001111000000000000100100000;
11'd379: out <= 32'b00000000100111000000000000000000;
11'd380: out <= 32'b00000001100001000000000000000000;
11'd381: out <= 32'b00000000000100000000000000001000;
11'd382: out <= 32'b00000001111000000000000100100000;
11'd383: out <= 32'b00000000000100000000000000001001;
11'd384: out <= 32'b00000001111000000000000100100000;
11'd385: out <= 32'b00000000010011000000000000000000;
11'd386: out <= 32'b00000000010010000000000000000000;
11'd387: out <= 32'b00000001011110100000000000000111;
11'd388: out <= 32'b00000001010000000000000110000110;
11'd389: out <= 32'b00000000010100000000000101111000;
11'd390: out <= 32'b00000000011100000010000100011001;
11'd391: out <= 32'b00000001100001000000000000000000;
11'd392: out <= 32'b00000001011101010000000001111110;
11'd393: out <= 32'b00000001010000000000000110001101;
11'd394: out <= 32'b00000000010001000000000000000000;
11'd395: out <= 32'b00000000011001000000000000000000;
11'd396: out <= 32'b00000000010100000000000101110011;
11'd397: out <= 32'b00000000011100000010000100011001;
11'd398: out <= 32'b00000000000100000000000000000000;
11'd399: out <= 32'b00000000011000000000000000000000;
11'd400: out <= 32'b00000001111000000000000000001001;
11'd401: out <= 32'b00000001111100000000000000000000;
11'd402: out <= 32'b00000000000110000000000000000000;
11'd403: out <= 32'b00000000000100000000000000000011;
11'd404: out <= 32'b00000001100101100000000000000000;
11'd405: out <= 32'b00000001111000000000000100100000;
11'd406: out <= 32'b00000000000100000000000000000100;
11'd407: out <= 32'b00000000000101000000000000000000;
11'd408: out <= 32'b00000001111000000000000100100000;
11'd409: out <= 32'b00000000000100000000000000000101;
11'd410: out <= 32'b00000000000101000000000000000000;
11'd411: out <= 32'b00000001111000000000000100100000;
11'd412: out <= 32'b00000000010011000000000000000000;
11'd413: out <= 32'b00000000010010000000000000000000;
11'd414: out <= 32'b00000001011110100000000000000010;
11'd415: out <= 32'b00000001010000000000000110100001;
11'd416: out <= 32'b00000000010100000000000110010011;
11'd417: out <= 32'b00000001111100000000000000000000;
11'd418: out <= 32'b00000000011100000010000000000010;
11'd419: out <= 32'b00000001100000000000000000000000;
11'd420: out <= 32'b00000001011100001111111111111111;
11'd421: out <= 32'b00000001001000000000000110100111;
11'd422: out <= 32'b00000000010100000000000110100010;
11'd423: out <= 32'b00000001111100000000000000000000;
11'd424: out <= 32'b00000001111000000000000000001001;
11'd425: out <= 32'b00000000011100000010000000000010;
11'd426: out <= 32'b00000000000100000000000000000000;
11'd427: out <= 32'b00000000011000000000000000000000;
11'd428: out <= 32'b00000000000100000000000011111101;
11'd429: out <= 32'b00000000000101000000000000000000;
11'd430: out <= 32'b00000001111000000000000100100000;
11'd431: out <= 32'b00000001111000000000000110100010;
11'd432: out <= 32'b00000001111100000000000000000000;
11'd433: out <= 32'b00000001111000000000000000001001;
11'd434: out <= 32'b00000000000101000000000000001000;
11'd435: out <= 32'b00000000011100000010000100010110;
11'd436: out <= 32'b00000000011001000000000000000000;
11'd437: out <= 32'b00000000011100000010000100010110;
11'd438: out <= 32'b00000001100001000000000000000000;
11'd439: out <= 32'b00000000000110000001101100000000;
11'd440: out <= 32'b00000001111000000000000101010110;
11'd441: out <= 32'b00000000011100000010000100010110;
11'd442: out <= 32'b00000001100001000000000000000000;
11'd443: out <= 32'b00000001011101010000000000011111;
11'd444: out <= 32'b00000001001000000000000111000000;
11'd445: out <= 32'b00000000010001000000000000000000;
11'd446: out <= 32'b00000000011001000000000000000000;
11'd447: out <= 32'b00000000010100000000000110110101;
11'd448: out <= 32'b00000001111100000000000000000000;
11'd449: out <= 32'b00000001111000000000000000010111;
11'd450: out <= 32'b00000000011100000001111111000010;
11'd451: out <= 32'b00000000000100000000000000000000;
11'd452: out <= 32'b00000000011000000000000000000000;
11'd453: out <= 32'b00000001100000000000000000000000;
11'd454: out <= 32'b00000001011100001111111111111111;
11'd455: out <= 32'b00000001001000000000000111001001;
11'd456: out <= 32'b00000000010100000000000111000101;
11'd457: out <= 32'b00000001111000000000000000100100;
11'd458: out <= 32'b00000001111100000000000000000000;
11'd459: out <= 32'b00000000110100000000000011111111;
11'd460: out <= 32'b00000001011100000000000011100000;
11'd461: out <= 32'b00000001001000000000000111011111;
11'd462: out <= 32'b00000001011100000000000000000000;
11'd463: out <= 32'b00000001001000000000001000100001;
11'd464: out <= 32'b00000001011100000000000011111111;
11'd465: out <= 32'b00000001001000000000001000100001;
11'd466: out <= 32'b00000001011100000000000011110000;
11'd467: out <= 32'b00000001001000000000000111100010;
11'd468: out <= 32'b00000000011100000010000100000011;
11'd469: out <= 32'b00000001100001000000000000000000;
11'd470: out <= 32'b00000000000110001111111111111111;
11'd471: out <= 32'b00000001011110010000000000000000;
11'd472: out <= 32'b00000001001000000000000111011010;
11'd473: out <= 32'b00000000010100000000001000100001;
11'd474: out <= 32'b00000000000101000000000000000000;
11'd475: out <= 32'b00000000011001000000000000000000;
11'd476: out <= 32'b00000001011100000000000001011001;
11'd477: out <= 32'b00000001001000000000000111101000;
11'd478: out <= 32'b00000000010100000000000111110010;
11'd479: out <= 32'b00000000011100000010000100000101;
11'd480: out <= 32'b00000000011000001111111111111111;
11'd481: out <= 32'b00000000010100000000000111100100;
11'd482: out <= 32'b00000000011100000010000100000101;
11'd483: out <= 32'b00000000011000000000000000000000;
11'd484: out <= 32'b00000000011100000010000100000011;
11'd485: out <= 32'b00000000011000001111111111111111;
11'd486: out <= 32'b00000000000100000000000000000000;
11'd487: out <= 32'b00000000010100000000001000011001;
11'd488: out <= 32'b00000000011100000010000100000100;
11'd489: out <= 32'b00000001100000000000000000000000;
11'd490: out <= 32'b00000000000101001111111111111111;
11'd491: out <= 32'b00000001011100010000000000000000;
11'd492: out <= 32'b00000001001000000000000111101111;
11'd493: out <= 32'b00000000011000001111111111111111;
11'd494: out <= 32'b00000000010100000000001000100001;
11'd495: out <= 32'b00000000000101000000000000000000;
11'd496: out <= 32'b00000000011001000000000000000000;
11'd497: out <= 32'b00000000010100000000001000100001;
11'd498: out <= 32'b00000000000101000000011111000000;
11'd499: out <= 32'b00000000000111000000000000000000;
11'd500: out <= 32'b00000000100101000000000000000000;
11'd501: out <= 32'b00000001100010000000000000000000;
11'd502: out <= 32'b00000000011100000010000100000000;
11'd503: out <= 32'b00000000011001000000000000000000;
11'd504: out <= 32'b00000000011100000010000100000001;
11'd505: out <= 32'b00000000011011000000000000000000;
11'd506: out <= 32'b00000000011100000010000100000100;
11'd507: out <= 32'b00000001100001000000000000000000;
11'd508: out <= 32'b00000001011101011111111111111111;
11'd509: out <= 32'b00000001001000000000001000000000;
11'd510: out <= 32'b00000000110110000000000011111111;
11'd511: out <= 32'b00000000010100000000001000000011;
11'd512: out <= 32'b00000000000111000000000000000111;
11'd513: out <= 32'b00000001000010110000000000000000;
11'd514: out <= 32'b00000001001110000000000000000000;
11'd515: out <= 32'b00000000011100000010000100000000;
11'd516: out <= 32'b00000001100001000000000000000000;
11'd517: out <= 32'b00000000011100000010000100000001;
11'd518: out <= 32'b00000001100011000000000000000000;
11'd519: out <= 32'b00000001011100100000000000000000;
11'd520: out <= 32'b00000001001000000000001000001111;
11'd521: out <= 32'b00000000000110000000000000111111;
11'd522: out <= 32'b00000001011110110000000000000000;
11'd523: out <= 32'b00000001001000000000001000001101;
11'd524: out <= 32'b00000000010100000000001000010001;
11'd525: out <= 32'b00000000000100000000000000000000;
11'd526: out <= 32'b00000000010100000000001000010100;
11'd527: out <= 32'b00000001100100110000000000000000;
11'd528: out <= 32'b00000000010100000000001000010100;
11'd529: out <= 32'b00000000010011000000000000000000;
11'd530: out <= 32'b00000000010001000000000000000000;
11'd531: out <= 32'b00000000010100000000000111110100;
11'd532: out <= 32'b00000000011100000010000100000100;
11'd533: out <= 32'b00000000000101000000000000000000;
11'd534: out <= 32'b00000000011001000000000000000000;
11'd535: out <= 32'b00000000010100000000001000011001;
11'd536: out <= 32'b00000000000100000000000000000000;
11'd537: out <= 32'b00000000000101000000000000000000;
11'd538: out <= 32'b00000001011100010000000000000000;
11'd539: out <= 32'b00000001001000000000001000100001;
11'd540: out <= 32'b00000000011100000001111111100001;
11'd541: out <= 32'b00000000011000000000000000000000;
11'd542: out <= 32'b00000000011100000010000100000110;
11'd543: out <= 32'b00000000011000001111111111111111;
11'd544: out <= 32'b00000000010100000000001000100100;
11'd545: out <= 32'b00000000011100000010000100000110;
11'd546: out <= 32'b00000000000101000000000000000000;
11'd547: out <= 32'b00000000011001000000000000000000;
11'd548: out <= 32'b00000001111000000000000000101101;
11'd549: out <= 32'b00000001111100000000000000000000;
11'd550: out <= 32'b00000001111000000000000000011010;
11'd551: out <= 32'b00000000011100000010000100010001;
11'd552: out <= 32'b00000001100000000000000000000000;
11'd553: out <= 32'b00000001011100001111111111111111;
11'd554: out <= 32'b00000001001000000000001000101110;
11'd555: out <= 32'b00000000000011000000000000000011;
11'd556: out <= 32'b00000000001000000000000000000000;
11'd557: out <= 32'b00000001111000000000000111001011;
11'd558: out <= 32'b00000001111000000000000000101101;
11'd559: out <= 32'b00000001111100000000000000000000;
11'd560: out <= 32'b00000000011100000010000100010010;
11'd561: out <= 32'b00000000011000000000000000000000;
11'd562: out <= 32'b00000000001101000000000000000000;
11'd563: out <= 32'b00000000001100000000000000000001;
11'd564: out <= 32'b00000001111100000000000000000000;
11'd565: out <= 32'b00000000011100000010000100010010;
11'd566: out <= 32'b00000001100001000000000000000000;
11'd567: out <= 32'b00000001011101011111111111111111;
11'd568: out <= 32'b00000001001000000000001000111010;
11'd569: out <= 32'b00000000010100000000001000110101;
11'd570: out <= 32'b00000000011000000000000000000000;
11'd571: out <= 32'b00000001111100000000000000000000;
11'd572: out <= 32'b00000001111000000000000000011010;
11'd573: out <= 32'b00000000000011000000000000000000;
11'd574: out <= 32'b00000000001000000000000000000000;
11'd575: out <= 32'b00000000011100000010000100010101;
11'd576: out <= 32'b00000000011000000000000000000000;
11'd577: out <= 32'b00000000011100000010000100010010;
11'd578: out <= 32'b00000000011000001111111111111111;
11'd579: out <= 32'b00000001111000000000000000101101;
11'd580: out <= 32'b00000001111100000000000000000000;
11'd581: out <= 32'b00000000000100000000000000000001;
11'd582: out <= 32'b00000000000101000000000000000000;
11'd583: out <= 32'b00000001111000000000001000110000;
11'd584: out <= 32'b00000001111000000000001000110101;
11'd585: out <= 32'b00000001111100000000000000000000;
11'd586: out <= 32'b00000000011100000010000100010001;
11'd587: out <= 32'b00000000011000001111111111111111;
11'd588: out <= 32'b00000001111100000000000000000000;
11'd589: out <= 32'b00000000011100000010000100010001;
11'd590: out <= 32'b00000000011000000000000000000000;
11'd591: out <= 32'b00000001111100000000000000000000;
11'd592: out <= 32'b00000001111000000000000000010111;
11'd593: out <= 32'b00000001111000000000001001001010;
11'd594: out <= 32'b00000001111000000000001001000101;
11'd595: out <= 32'b00000001111000000000000000100100;
11'd596: out <= 32'b00000001111100000000000000000000;
11'd597: out <= 32'b00000001111000000000000000010111;
11'd598: out <= 32'b00000000000100000000000000000010;
11'd599: out <= 32'b00000000011100000010000100011000;
11'd600: out <= 32'b00000001100001000000000000000000;
11'd601: out <= 32'b00000001111000000000001000110000;
11'd602: out <= 32'b00000000000111000000000000000000;
11'd603: out <= 32'b00000000000110000000000000000000;
11'd604: out <= 32'b00000000000100000000000000000011;
11'd605: out <= 32'b00000000000101000000000000000000;
11'd606: out <= 32'b00000001111000000000001000110000;
11'd607: out <= 32'b00000001111000000000001000110101;
11'd608: out <= 32'b00000000011100000010000100010100;
11'd609: out <= 32'b00000000011000000000000000000000;
11'd610: out <= 32'b00000000000100000000000000000101;
11'd611: out <= 32'b00000000000101000000000000000000;
11'd612: out <= 32'b00000001111000000000001000110000;
11'd613: out <= 32'b00000001111000000000001000110101;
11'd614: out <= 32'b00000000000111000000000000000000;
11'd615: out <= 32'b00000000000100000000000000000111;
11'd616: out <= 32'b00000000000101000000000000000000;
11'd617: out <= 32'b00000001111000000000001000110000;
11'd618: out <= 32'b00000000011100000010000100010100;
11'd619: out <= 32'b00000001100000000000000000000000;
11'd620: out <= 32'b00000001011100001111111111111111;
11'd621: out <= 32'b00000001001000000000001001111010;
11'd622: out <= 32'b00000000011000001111111111111111;
11'd623: out <= 32'b00000000011100000010000100010101;
11'd624: out <= 32'b00000001100000000000000000000000;
11'd625: out <= 32'b00000000000101000000000000000111;
11'd626: out <= 32'b00000000111100010000000000000000;
11'd627: out <= 32'b00000001001100000000000000000000;
11'd628: out <= 32'b00000000011100000010000100010011;
11'd629: out <= 32'b00000001100001000000000000000000;
11'd630: out <= 32'b00000000100101000000000000000000;
11'd631: out <= 32'b00000001100001000000000000000000;
11'd632: out <= 32'b00000000011000000000000000000000;
11'd633: out <= 32'b00000000010100000000001010001000;
11'd634: out <= 32'b00000000000100000000000000000000;
11'd635: out <= 32'b00000000011000000000000000000000;
11'd636: out <= 32'b00000000011100000010000100010101;
11'd637: out <= 32'b00000001100000000000000000000000;
11'd638: out <= 32'b00000000011100000010000100010011;
11'd639: out <= 32'b00000001100001000000000000000000;
11'd640: out <= 32'b00000000100101000000000000000000;
11'd641: out <= 32'b00000001100001000000000000000000;
11'd642: out <= 32'b00000000111000010000000000000000;
11'd643: out <= 32'b00000000011000000000000000000000;
11'd644: out <= 32'b00000000011100000010000100010011;
11'd645: out <= 32'b00000001100000000000000000000000;
11'd646: out <= 32'b00000000010000000000000000000000;
11'd647: out <= 32'b00000000011000000000000000000000;
11'd648: out <= 32'b00000001011111110000000000000111;
11'd649: out <= 32'b00000001001000000000001010001100;
11'd650: out <= 32'b00000000010011000000000000000000;
11'd651: out <= 32'b00000000010100000000001001100111;
11'd652: out <= 32'b00000001011110100000000000111111;
11'd653: out <= 32'b00000001001000000000001010010000;
11'd654: out <= 32'b00000000010010000000000000000000;
11'd655: out <= 32'b00000000010100000000001001100010;
11'd656: out <= 32'b00000001111000000000001001001101;
11'd657: out <= 32'b00000001111000000000000000100100;
11'd658: out <= 32'b00000001111100000000000000000000;
11'd659: out <= 32'b00000000011100000010000100010011;
11'd660: out <= 32'b00000000011000000001000000000000;
11'd661: out <= 32'b00000000011100000010000100011000;
11'd662: out <= 32'b00000000000100000000000000000000;
11'd663: out <= 32'b00000000011000000000000000000000;
11'd664: out <= 32'b00000001111000000000001001010101;
11'd665: out <= 32'b00000000011100000010000100010011;
11'd666: out <= 32'b00000001100000000000000000000000;
11'd667: out <= 32'b00000001011100000001001111111111;
11'd668: out <= 32'b00000001010000000000001010100011;
11'd669: out <= 32'b00000001001000000000001010100011;
11'd670: out <= 32'b00000000011100000010000100011000;
11'd671: out <= 32'b00000001100000000000000000000000;
11'd672: out <= 32'b00000000010000000000000000000000;
11'd673: out <= 32'b00000000011000000000000000000000;
11'd674: out <= 32'b00000000010100000000001010011000;
11'd675: out <= 32'b00000000011100000001000011111111;
11'd676: out <= 32'b00000001100000000000000000000000;
11'd677: out <= 32'b00000000011100000001111111100001;
11'd678: out <= 32'b00000000011000000000000000000000;
11'd679: out <= 32'b00000001111100000000000000000000;
11'd680: out <= 32'b00000001111000000000000000001001;
11'd681: out <= 32'b00000000011100000001111110100101;
11'd682: out <= 32'b00000000000111000000000000000000;
11'd683: out <= 32'b00000000011011000000000000000000;
11'd684: out <= 32'b00000000000110000001111110101000;
11'd685: out <= 32'b00000000100110000000000000000000;
11'd686: out <= 32'b00000000011000000000000000000000;
11'd687: out <= 32'b00000000010010000000000000000000;
11'd688: out <= 32'b00000001011110100001111110101101;
11'd689: out <= 32'b00000001010100000000001010101101;
11'd690: out <= 32'b00000000011100000001111110101101;
11'd691: out <= 32'b00000000011000000000000000001111;
11'd692: out <= 32'b00000000011100000001111110100100;
11'd693: out <= 32'b00000001100000000000000000000000;
11'd694: out <= 32'b00000001100110000000000000000000;
11'd695: out <= 32'b00000000110100001000000000000000;
11'd696: out <= 32'b00000000000101000000000000000111;
11'd697: out <= 32'b00000001000000010000000000000000;
11'd698: out <= 32'b00000001001100000000000000000000;
11'd699: out <= 32'b00000000000101000000000000000110;
11'd700: out <= 32'b00000001000000010000000000000000;
11'd701: out <= 32'b00000001001100000000000000000000;
11'd702: out <= 32'b00000001100111000000000000000000;
11'd703: out <= 32'b00000000000101000000000000000000;
11'd704: out <= 32'b00000000111110010000000000000000;
11'd705: out <= 32'b00000001001110000000000000000000;
11'd706: out <= 32'b00000000110110001111111111111111;
11'd707: out <= 32'b00000000011010000000000000000000;
11'd708: out <= 32'b00000000011100000001111110101110;
11'd709: out <= 32'b00000000011000000001111110101101;
11'd710: out <= 32'b00000000011100000001111110101110;
11'd711: out <= 32'b00000001100000000000000000000000;
11'd712: out <= 32'b00000001011000000000000000000000;
11'd713: out <= 32'b00000000011000000000000000000000;
11'd714: out <= 32'b00000000100100000000000000000000;
11'd715: out <= 32'b00000001100000000000000000000000;
11'd716: out <= 32'b00000001011100000000000000000101;
11'd717: out <= 32'b00000001001000000000001011010000;
11'd718: out <= 32'b00000001010000000000001011010000;
11'd719: out <= 32'b00000000010100000000001011010001;
11'd720: out <= 32'b00000000101100000000000000000011;
11'd721: out <= 32'b00000001100110000000000000000000;
11'd722: out <= 32'b00000000110110000000000000001000;
11'd723: out <= 32'b00000000000101000000000000000010;
11'd724: out <= 32'b00000001000010010000000000000000;
11'd725: out <= 32'b00000001001110000000000000000000;
11'd726: out <= 32'b00000000000101000000000000000000;
11'd727: out <= 32'b00000000111100010000000000000000;
11'd728: out <= 32'b00000001001100000000000000000000;
11'd729: out <= 32'b00000000101100110000000000000000;
11'd730: out <= 32'b00000000110100000000000000001111;
11'd731: out <= 32'b00000001100111100000000000000000;
11'd732: out <= 32'b00000000011000000000000000000000;
11'd733: out <= 32'b00000000011100000001111110101110;
11'd734: out <= 32'b00000001100000000000000000000000;
11'd735: out <= 32'b00000001011100000001111110101001;
11'd736: out <= 32'b00000001010000000000001011000110;
11'd737: out <= 32'b00000000011100000001111110101000;
11'd738: out <= 32'b00000001100000000000000000000000;
11'd739: out <= 32'b00000001011100000000000000000101;
11'd740: out <= 32'b00000001001000000000001011100111;
11'd741: out <= 32'b00000001010000000000001011100111;
11'd742: out <= 32'b00000000010100000000001011101000;
11'd743: out <= 32'b00000000101100000000000000000011;
11'd744: out <= 32'b00000001100110000000000000000000;
11'd745: out <= 32'b00000000000101000000000000000000;
11'd746: out <= 32'b00000000111100010000000000000000;
11'd747: out <= 32'b00000001001100000000000000000000;
11'd748: out <= 32'b00000000101100110000000000000000;
11'd749: out <= 32'b00000000110100000000000000001111;
11'd750: out <= 32'b00000000011000000000000000000000;
11'd751: out <= 32'b00000000011100000001111110100101;
11'd752: out <= 32'b00000001100000000000000000000000;
11'd753: out <= 32'b00000001011100000000000000001110;
11'd754: out <= 32'b00000001010000000000001011110110;
11'd755: out <= 32'b00000000010000000000000000000000;
11'd756: out <= 32'b00000000011000000000000000000000;
11'd757: out <= 32'b00000000010100000000001010110100;
11'd758: out <= 32'b00000000000100000001111110101000;
11'd759: out <= 32'b00000000100100000000000000000000;
11'd760: out <= 32'b00000001100011000000000000000000;
11'd761: out <= 32'b00000000010011000000000000000000;
11'd762: out <= 32'b00000000011011000000000000000000;
11'd763: out <= 32'b00000000010000000000000000000000;
11'd764: out <= 32'b00000001011100000001111110101101;
11'd765: out <= 32'b00000001001000000000001011111111;
11'd766: out <= 32'b00000000010100000000001011110111;
11'd767: out <= 32'b00000001111100000000000000000000;
11'd768: out <= 32'b00000000011100000001111110100100;
11'd769: out <= 32'b00000001100000000000000000000000;
11'd770: out <= 32'b00000001011100000000000000000000;
11'd771: out <= 32'b00000001010100000000001100000101;
11'd772: out <= 32'b00000000010100000000001100001000;
11'd773: out <= 32'b00000000011100000001111110110001;
11'd774: out <= 32'b00000000011000000000000000001011;
11'd775: out <= 32'b00000000010100000000001100001100;
11'd776: out <= 32'b00000000011100000001111110110001;
11'd777: out <= 32'b00000000000101000000000000000000;
11'd778: out <= 32'b00000000011001000000000000000000;
11'd779: out <= 32'b00000000010100000000001100001100;
11'd780: out <= 32'b00000000011100000001111110100100;
11'd781: out <= 32'b00000001111000000000000001110000;
11'd782: out <= 32'b00000000011000000000000000000000;
11'd783: out <= 32'b00000001111000000000001010101000;
11'd784: out <= 32'b00000000000101000001111110101000;
11'd785: out <= 32'b00000000000110000001111110110010;
11'd786: out <= 32'b00000000100101000000000000000000;
11'd787: out <= 32'b00000001100011000000000000000000;
11'd788: out <= 32'b00000000100110000000000000000000;
11'd789: out <= 32'b00000000011011000000000000000000;
11'd790: out <= 32'b00000000010001000000000000000000;
11'd791: out <= 32'b00000000010010000000000000000000;
11'd792: out <= 32'b00000001011101010001111110101101;
11'd793: out <= 32'b00000001001000000000001100011011;
11'd794: out <= 32'b00000000010100000000001100010010;
11'd795: out <= 32'b00000000011100000001111110110111;
11'd796: out <= 32'b00000000011000000000000000001111;
11'd797: out <= 32'b00000001111000000000001100011111;
11'd798: out <= 32'b00000001111100000000000000000000;
11'd799: out <= 32'b00000000011100000001111110110011;
11'd800: out <= 32'b00000001100000000000000000000000;
11'd801: out <= 32'b00000001011100000000000000111010;
11'd802: out <= 32'b00000001001000000000001100111011;
11'd803: out <= 32'b00000001011100000000000000001111;
11'd804: out <= 32'b00000001001000000000001100111011;
11'd805: out <= 32'b00000000011100000001111110110010;
11'd806: out <= 32'b00000001100000000000000000000000;
11'd807: out <= 32'b00000001011100000000000000000000;
11'd808: out <= 32'b00000001001000000000001100101100;
11'd809: out <= 32'b00000001011100000000000000000001;
11'd810: out <= 32'b00000001001000000000001100101100;
11'd811: out <= 32'b00000000010100000000001100111011;
11'd812: out <= 32'b00000000000100000001111110110011;
11'd813: out <= 32'b00000000100100000000000000000000;
11'd814: out <= 32'b00000001100011000000000000000000;
11'd815: out <= 32'b00000001011000000000000000000000;
11'd816: out <= 32'b00000000100100000000000000000000;
11'd817: out <= 32'b00000000011011000000000000000000;
11'd818: out <= 32'b00000000010000000000000000000000;
11'd819: out <= 32'b00000000010000000000000000000000;
11'd820: out <= 32'b00000001011100000001111110111011;
11'd821: out <= 32'b00000001001000000000001100110111;
11'd822: out <= 32'b00000000010100000000001100101101;
11'd823: out <= 32'b00000000011100000001111110111010;
11'd824: out <= 32'b00000000000111000000000000000000;
11'd825: out <= 32'b00000000011011000000000000000000;
11'd826: out <= 32'b00000000010100000000001100011111;
11'd827: out <= 32'b00000001111100000000000000000000;
11'd828: out <= 32'b00000000000100000000000000001010;
11'd829: out <= 32'b00000000011100000001111111000000;
11'd830: out <= 32'b00000001100001000000000000000000;
11'd831: out <= 32'b00000000000110000000000000000010;
11'd832: out <= 32'b00000000111101100000000000000000;
11'd833: out <= 32'b00000001001101000000000000000000;
11'd834: out <= 32'b00000001111000000000000100100000;
11'd835: out <= 32'b00000000000100000000000000001011;
11'd836: out <= 32'b00000000011100000001111111000001;
11'd837: out <= 32'b00000001100001000000000000000000;
11'd838: out <= 32'b00000000000110000000000000000010;
11'd839: out <= 32'b00000000111101100000000000000000;
11'd840: out <= 32'b00000001001101000000000000000000;
11'd841: out <= 32'b00000001111000000000000100100000;
11'd842: out <= 32'b00000000000100000000000000001100;
11'd843: out <= 32'b00000001111100000000000000000000;
11'd844: out <= 32'b00000001111000000000000000001001;
11'd845: out <= 32'b00000000000111000000000000000000;
11'd846: out <= 32'b00000001111000000000001100111100;
11'd847: out <= 32'b00000000011100000001111111000011;
11'd848: out <= 32'b00000001100001000000000000000000;
11'd849: out <= 32'b00000001100110010000000000000000;
11'd850: out <= 32'b00000000010010000000000000000000;
11'd851: out <= 32'b00000000011010000000000000000000;
11'd852: out <= 32'b00000000100101000000000000000000;
11'd853: out <= 32'b00000001100001000000000000000000;
11'd854: out <= 32'b00000000011100000010000100010110;
11'd855: out <= 32'b00000001100000000000000000000000;
11'd856: out <= 32'b00000001011100001111111111111111;
11'd857: out <= 32'b00000001001000000000001101011100;
11'd858: out <= 32'b00000000110101000000000011111111;
11'd859: out <= 32'b00000000010100000000001101011111;
11'd860: out <= 32'b00000000000100000000000000000111;
11'd861: out <= 32'b00000001000001000000000000000000;
11'd862: out <= 32'b00000001001101000000000000000000;
11'd863: out <= 32'b00000000000100000000000000001100;
11'd864: out <= 32'b00000001011101010000000000010000;
11'd865: out <= 32'b00000001001000000000001101101011;
11'd866: out <= 32'b00000001011101010000000000001111;
11'd867: out <= 32'b00000001001000000000001101111010;
11'd868: out <= 32'b00000001111000000000000100100000;
11'd869: out <= 32'b00000001111000000000000001101011;
11'd870: out <= 32'b00000000011100000001111111000000;
11'd871: out <= 32'b00000001100001000000000000000000;
11'd872: out <= 32'b00000001011101010000000000100100;
11'd873: out <= 32'b00000001010000000000001101101011;
11'd874: out <= 32'b00000000010100000000001101110001;
11'd875: out <= 32'b00000000011100000001111111000000;
11'd876: out <= 32'b00000000011000000000000000000100;
11'd877: out <= 32'b00000000011100000001111111000001;
11'd878: out <= 32'b00000001100001000000000000000000;
11'd879: out <= 32'b00000000010001000000000000000000;
11'd880: out <= 32'b00000000011001000000000000000000;
11'd881: out <= 32'b00000000011100000001111111000000;
11'd882: out <= 32'b00000001100001000000000000000000;
11'd883: out <= 32'b00000000010001000000000000000000;
11'd884: out <= 32'b00000000011001000000000000000000;
11'd885: out <= 32'b00000000010011000000000000000000;
11'd886: out <= 32'b00000001011111110000000000111010;
11'd887: out <= 32'b00000001001000000000001101111010;
11'd888: out <= 32'b00000001010000000000001101111010;
11'd889: out <= 32'b00000000010100000000001101001110;
11'd890: out <= 32'b00000001111100000000000000000000;
11'd891: out <= 32'b00000001111000000000000000010111;
11'd892: out <= 32'b00000001111000000000001101001100;
11'd893: out <= 32'b00000001111000000000000000100100;
11'd894: out <= 32'b00000001111100000000000000000000;
11'd895: out <= 32'b00000001111000000000000000010111;
11'd896: out <= 32'b00000001111000000000001100000000;
11'd897: out <= 32'b00000000011100000001111111000011;
11'd898: out <= 32'b00000000000101000001111110110001;
11'd899: out <= 32'b00000000011001000000000000000000;
11'd900: out <= 32'b00000001111000000000001101001100;
11'd901: out <= 32'b00000001111000000000000000100100;
11'd902: out <= 32'b00000001111100000000000000000000;
11'd903: out <= 32'b00000001111000000000000000010111;
11'd904: out <= 32'b00000000011100000010000100000101;
11'd905: out <= 32'b00000001100000000000000000000000;
11'd906: out <= 32'b00000001011100001111111111111111;
11'd907: out <= 32'b00000001001000000000001110001101;
11'd908: out <= 32'b00000000010100000000001110001000;
11'd909: out <= 32'b00000001111000000000000000100100;
11'd910: out <= 32'b00000001111100000000000000000000;
11'd911: out <= 32'b00000000011100000010000100000101;
11'd912: out <= 32'b00000000011000000000000000000000;
11'd913: out <= 32'b00000001111100000000000000000000;
11'd914: out <= 32'b00000001111000000000000000010111;
11'd915: out <= 32'b00000001111000000000001110001111;
11'd916: out <= 32'b00000001111000000000000000100100;
11'd917: out <= 32'b00000001111100000000000000000000;
11'd918: out <= 32'b00000001111000000000000000010111;
11'd919: out <= 32'b00000001111000000000001110001111;
11'd920: out <= 32'b00000001111000000000000000100100;
11'd921: out <= 32'b00000001111100000000000000000000;
11'd922: out <= 32'b11010111001010110100010100100101;
11'd923: out <= 32'b00000001001011110100111100011101;
11'd924: out <= 32'b11010111110110111011010001011111;
11'd925: out <= 32'b11001000001101110100110000111111;
11'd926: out <= 32'b00010010111010010111100100001110;
11'd927: out <= 32'b10100000011011010001011100111010;
11'd928: out <= 32'b01000001011000011011110000110010;
11'd929: out <= 32'b01100010001100110000100110111000;
11'd930: out <= 32'b11101110101110010000011001100110;
11'd931: out <= 32'b10001100010000111000011000001000;
11'd932: out <= 32'b10100011100110010111100111001001;
11'd933: out <= 32'b01101000011101011100110000100110;
11'd934: out <= 32'b10100101100111110110101100111010;
11'd935: out <= 32'b11000110101011000110000010000100;
11'd936: out <= 32'b11010010010001010011011110010000;
11'd937: out <= 32'b10110111101011011101000111101010;
11'd938: out <= 32'b00011011101101010010101010000111;
11'd939: out <= 32'b10101011110100101010011000101010;
11'd940: out <= 32'b10101001101001011010011101111110;
11'd941: out <= 32'b00101111110101000100100000111000;
11'd942: out <= 32'b00001011110010001011001001000010;
11'd943: out <= 32'b11101110100001100010011101101011;
11'd944: out <= 32'b01100000110011001011010101111111;
11'd945: out <= 32'b11011110000100000001100101010001;
11'd946: out <= 32'b10100010001000000000010000011011;
11'd947: out <= 32'b01010101001100000100100101000100;
11'd948: out <= 32'b00001111100011010101010000110100;
11'd949: out <= 32'b01100001000101110100000111110101;
11'd950: out <= 32'b11100000111100010001000010011010;
11'd951: out <= 32'b00101000011010001001100010100011;
11'd952: out <= 32'b10011111000010011110100010011101;
11'd953: out <= 32'b00001111000001000100010001001011;
11'd954: out <= 32'b01000010001111101000011000110010;
11'd955: out <= 32'b01101111101000000100111000100101;
11'd956: out <= 32'b01001011011101000010100000000001;
11'd957: out <= 32'b00000001100010000000111001100011;
11'd958: out <= 32'b10101001110010010001011111001110;
11'd959: out <= 32'b11110111101100111000010101011101;
11'd960: out <= 32'b00110110110111011100010010001010;
11'd961: out <= 32'b00011000000110101101001010011010;
11'd962: out <= 32'b01101011011110001000111110110000;
11'd963: out <= 32'b11001111101101100011010000110010;
11'd964: out <= 32'b00110000001001010000110011111100;
11'd965: out <= 32'b11110010000100011000110010101001;
11'd966: out <= 32'b00101000001100011000001100111001;
11'd967: out <= 32'b00111100010100010101111011011000;
11'd968: out <= 32'b01100011101111011001100111100011;
11'd969: out <= 32'b01100111011000011100010111011010;
11'd970: out <= 32'b00001100011001100111111000110101;
11'd971: out <= 32'b10000001011100011011000011111111;
11'd972: out <= 32'b11110000000101000011000100101001;
11'd973: out <= 32'b10100001000101001101011010010000;
11'd974: out <= 32'b01100100011001000000100010010010;
11'd975: out <= 32'b01000111110110001010100011110011;
11'd976: out <= 32'b01001001101000001110111011010001;
11'd977: out <= 32'b00000011010000010001011000110111;
11'd978: out <= 32'b10001001110010100011100111101111;
11'd979: out <= 32'b10111011100110001001101010001001;
11'd980: out <= 32'b00011010111110100000111101100110;
11'd981: out <= 32'b01101010111111100110000101010111;
11'd982: out <= 32'b01000000111010001111010011010011;
11'd983: out <= 32'b00111111100001101101010001111111;
11'd984: out <= 32'b00100000001010000011000100100001;
11'd985: out <= 32'b00100100001000010011001100101011;
11'd986: out <= 32'b00000000001100010010001100100100;
11'd987: out <= 32'b00100111001110000010001000110001;
11'd988: out <= 32'b00101111001010000010100000000000;
11'd989: out <= 32'b00110101001100110000000000101101;
11'd990: out <= 32'b00000010001001100000000100100100;
11'd991: out <= 32'b10100001000010110000111100001111;
11'd992: out <= 32'b00000000010001010000000000000000;
11'd993: out <= 32'b00011110000111100000000000010110;
11'd994: out <= 32'b00000000001001010010011000100110;
11'd995: out <= 32'b00110110001101100000000000101110;
11'd996: out <= 32'b00000000001111100011110100111101;
11'd997: out <= 32'b01001110010011100000000001000110;
11'd998: out <= 32'b00111110011111000101010101111001;
11'd999: out <= 32'b00000000011001100000000001001010;
11'd1000: out <= 32'b00000000011101010000000001011010;
11'd1001: out <= 32'b00000000011010110000000001110010;
11'd1002: out <= 32'b00010001000100010000000001110100;
11'd1003: out <= 32'b00010100000101000001010000101001;
11'd1004: out <= 32'b01000101000000000001001000010010;
11'd1005: out <= 32'b01000110000000000101001001010010;
11'd1006: out <= 32'b00101110000000000000000001010101;
11'd1007: out <= 32'b01001010000000000010010100000000;
11'd1008: out <= 32'b00110010001100100001110000011100;
11'd1009: out <= 32'b00100011001000110010000100100001;
11'd1010: out <= 32'b00101011001010110010010000100100;
11'd1011: out <= 32'b00110011001100110011010000110100;
11'd1012: out <= 32'b00111011001110110100001101000011;
11'd1013: out <= 32'b01001011010010110100001001000010;
11'd1014: out <= 32'b00110001001100010011101000111010;
11'd1015: out <= 32'b01001101010011010100010001000100;
11'd1016: out <= 32'b00101101001011010001010100010101;
11'd1017: out <= 32'b00101100001011000001101100011011;
11'd1018: out <= 32'b00101010001010100011110000111100;
11'd1019: out <= 32'b00100010001000100001110100011101;
11'd1020: out <= 32'b00011010000110100011010100110101;
11'd1021: out <= 32'b00000000010000010000000001001001;
11'd1022: out <= 32'b00000000010011000100110000000000;
11'd1023: out <= 32'b00010110000000000001111100011111;

default: out <= 0;
endcase
endmodule

module ROM2(
       input clk,
       input[7:0] addr,
       output reg[31:0] out
);

reg[31:0] memory[255:0];

initial begin
	memory[0] = 32'b00000000000000000000000000000000;
	memory[1] = 32'b00000000000000000000000000000000;
	memory[2] = 32'b00000000000000000000000000000000;
	memory[3] = 32'b00000000000000000000000000000000;
	memory[4] = 32'b00111100001111000000111111110000;
	memory[5] = 32'b00111111001111000011110011111100;
	memory[6] = 32'b00111100001111000011110000111100;
	memory[7] = 32'b00000000000000000000111111110000;
	memory[8] = 32'b00000011110000000000001111000000;
	memory[9] = 32'b00000011110000000000111111000000;
	memory[10] = 32'b00000011110000000000001111000000;
	memory[11] = 32'b00000000000000000011111111111100;
	memory[12] = 32'b00111100001111000000111111110000;
	memory[13] = 32'b00000000111100000000000000111100;
	memory[14] = 32'b00111100000000000000111100000000;
	memory[15] = 32'b00000000000000000011111111111100;
	memory[16] = 32'b00111100001111000000111111110000;
	memory[17] = 32'b00000011111100000000000000111100;
	memory[18] = 32'b00111100001111000000000000111100;
	memory[19] = 32'b00000000000000000000111111110000;
	memory[20] = 32'b00000000111111000000000000111100;
	memory[21] = 32'b00111100001111000000001111111100;
	memory[22] = 32'b00000000001111000011111111111111;
	memory[23] = 32'b00000000000000000000000000111100;
	memory[24] = 32'b00111100000000000011111111111100;
	memory[25] = 32'b00000000001111000011111111110000;
	memory[26] = 32'b00111100001111000000000000111100;
	memory[27] = 32'b00000000000000000000111111110000;
	memory[28] = 32'b00111100001111000000111111110000;
	memory[29] = 32'b00111111111100000011110000000000;
	memory[30] = 32'b00111100001111000011110000111100;
	memory[31] = 32'b00000000000000000000111111110000;
	memory[32] = 32'b00111100001111000011111111111100;
	memory[33] = 32'b00000011110000000000000011110000;
	memory[34] = 32'b00000011110000000000001111000000;
	memory[35] = 32'b00000000000000000000001111000000;
	memory[36] = 32'b00111100001111000000111111110000;
	memory[37] = 32'b00001111111100000011110000111100;
	memory[38] = 32'b00111100001111000011110000111100;
	memory[39] = 32'b00000000000000000000111111110000;
	memory[40] = 32'b00111100001111000000111111110000;
	memory[41] = 32'b00001111111111000011110000111100;
	memory[42] = 32'b00111100001111000000000000111100;
	memory[43] = 32'b00000000000000000000111111110000;
	memory[44] = 32'b00000000000000000000000000000000;
	memory[45] = 32'b00111111111111000000000000000000;
	memory[46] = 32'b00000000000000000000000000000000;
	memory[47] = 32'b00000000000000000000000000000000;
	memory[48] = 32'b00000011110000000000000000000000;
	memory[49] = 32'b00111111111111000000001111000000;
	memory[50] = 32'b00000011110000000000001111000000;
	memory[51] = 32'b00000000000000000000000000000000;
	memory[52] = 32'b00111100001111000000000000000000;
	memory[53] = 32'b11111111111111110000111111110000;
	memory[54] = 32'b00111100001111000000111111110000;
	memory[55] = 32'b00000000000000000000000000000000;
	memory[56] = 32'b00000000000011110000000000000000;
	memory[57] = 32'b00000000111100000000000000111100;
	memory[58] = 32'b00001111000000000000001111000000;
	memory[59] = 32'b00000000000000000011110000000000;
	memory[60] = 32'b11110000111100001111000011110000;
	memory[61] = 32'b00001111000011110000111100001111;
	memory[62] = 32'b11110000111100001111000011110000;
	memory[63] = 32'b00001111000011110000111100001111;
	memory[64] = 32'b11111111111111111111111111111111;
	memory[65] = 32'b11111111111111111111111111111111;
	memory[66] = 32'b11111111111111111111111111111111;
	memory[67] = 32'b11111111111111111111111111111111;
	memory[68] = 32'b11111111111111111111111111111111;
	memory[69] = 32'b11111111111111111111111111111111;
	memory[70] = 32'b00000000000000000000000000000000;
	memory[71] = 32'b00000000000000000000000000000000;
	memory[72] = 32'b00000000000000000000000000000000;
	memory[73] = 32'b00000000000000000000000000000000;
	memory[74] = 32'b11111111111111111111111111111111;
	memory[75] = 32'b11111111111111111111111111111111;
	memory[76] = 32'b11111111000000001111111100000000;
	memory[77] = 32'b11111111000000001111111100000000;
	memory[78] = 32'b11111111000000001111111100000000;
	memory[79] = 32'b11111111000000001111111100000000;
	memory[80] = 32'b00000000111111110000000011111111;
	memory[81] = 32'b00000000111111110000000011111111;
	memory[82] = 32'b00000000111111110000000011111111;
	memory[83] = 32'b00000000111111110000000011111111;
	memory[84] = 32'b11111100000011111111000000000011;
	memory[85] = 32'b00001111111111000011111100111111;
	memory[86] = 32'b00111111111111000000111111110000;
	memory[87] = 32'b11110000000011111111110000111111;
	memory[88] = 32'b00000000000000000000000000000000;
	memory[89] = 32'b00000000000000000000000000000000;
	memory[90] = 32'b00000000000000000000000000000000;
	memory[91] = 32'b11111111111111110000000000000000;
	memory[92] = 32'b00001111111100000000000000000000;
	memory[93] = 32'b00111111111111000011111111111100;
	memory[94] = 32'b00111111111111000011111111111100;
	memory[95] = 32'b00000000000000000000111111110000;
	memory[96] = 32'b00000011111100000000000011000000;
	memory[97] = 32'b00111111111111110000111111111100;
	memory[98] = 32'b00000011111100000000111111111100;
	memory[99] = 32'b00000000000000000000000011000000;
	memory[100] = 32'b00000011110000000011111100000000;
	memory[101] = 32'b00000000001111000000000011110000;
	memory[102] = 32'b00000011110000000000000011110000;
	memory[103] = 32'b00000000000000000011111100000000;
	memory[104] = 32'b00111100001111000011110000111100;
	memory[105] = 32'b00000000000000000011110000111100;
	memory[106] = 32'b00000000000000000000000000000000;
	memory[107] = 32'b00000000000000000000000000000000;
	memory[108] = 32'b00000011110000000000000011111100;
	memory[109] = 32'b00111100000000000000111100000000;
	memory[110] = 32'b00000011110000000000111100000000;
	memory[111] = 32'b00000000000000000000000011111100;
	memory[112] = 32'b00000000000000000000000000000000;
	memory[113] = 32'b00000000000000000011111111111100;
	memory[114] = 32'b00000000000000000011111111111100;
	memory[115] = 32'b00000000000000000000000000000000;
	memory[116] = 32'b00111100001111000011110000001100;
	memory[117] = 32'b00000011110000000000000011110000;
	memory[118] = 32'b00111100001111000000111100000000;
	memory[119] = 32'b00000000000000000011000000111100;
	memory[120] = 32'b00001111111111000000001111000000;
	memory[121] = 32'b00001111111100000011110000000000;
	memory[122] = 32'b00111111111100000000000000111100;
	memory[123] = 32'b00000000000000000000001111000000;
	memory[124] = 32'b00111100001111000000111111110000;
	memory[125] = 32'b00000000111100000000000000111100;
	memory[126] = 32'b00000000000000000000001111000000;
	memory[127] = 32'b00000000000000000000001111000000;
	memory[128] = 32'b00001111111100000000001111000000;
	memory[129] = 32'b00111111111111000011110000111100;
	memory[130] = 32'b00111100001111000011110000111100;
	memory[131] = 32'b00000000000000000011110000111100;
	memory[132] = 32'b00111100001111000011111111110000;
	memory[133] = 32'b00111111111100000011110000111100;
	memory[134] = 32'b00111100001111000011110000111100;
	memory[135] = 32'b00000000000000000011111111110000;
	memory[136] = 32'b00111100001111000000111111110000;
	memory[137] = 32'b00111100000000000011110000000000;
	memory[138] = 32'b00111100001111000011110000000000;
	memory[139] = 32'b00000000000000000000111111110000;
	memory[140] = 32'b00111100111100000011111111000000;
	memory[141] = 32'b00111100001111000011110000111100;
	memory[142] = 32'b00111100111100000011110000111100;
	memory[143] = 32'b00000000000000000011111111000000;
	memory[144] = 32'b00111100000000000011111111111100;
	memory[145] = 32'b00111111110000000011110000000000;
	memory[146] = 32'b00111100000000000011110000000000;
	memory[147] = 32'b00000000000000000011111111111100;
	memory[148] = 32'b00111100000000000011111111111100;
	memory[149] = 32'b00111111110000000011110000000000;
	memory[150] = 32'b00111100000000000011110000000000;
	memory[151] = 32'b00000000000000000011110000000000;
	memory[152] = 32'b00111100001111000000111111110000;
	memory[153] = 32'b00111100111111000011110000000000;
	memory[154] = 32'b00111100001111000011110000111100;
	memory[155] = 32'b00000000000000000000111111110000;
	memory[156] = 32'b00111100001111000011110000111100;
	memory[157] = 32'b00111111111111000011110000111100;
	memory[158] = 32'b00111100001111000011110000111100;
	memory[159] = 32'b00000000000000000011110000111100;
	memory[160] = 32'b00000011110000000000111111110000;
	memory[161] = 32'b00000011110000000000001111000000;
	memory[162] = 32'b00000011110000000000001111000000;
	memory[163] = 32'b00000000000000000000111111110000;
	memory[164] = 32'b00000000111100000000001111111100;
	memory[165] = 32'b00000000111100000000000011110000;
	memory[166] = 32'b00111100111100000000000011110000;
	memory[167] = 32'b00000000000000000000111111000000;
	memory[168] = 32'b00111100111100000011110000111100;
	memory[169] = 32'b00111111000000000011111111000000;
	memory[170] = 32'b00111100111100000011111111000000;
	memory[171] = 32'b00000000000000000011110000111100;
	memory[172] = 32'b00111100000000000011110000000000;
	memory[173] = 32'b00111100000000000011110000000000;
	memory[174] = 32'b00111100000000000011110000000000;
	memory[175] = 32'b00000000000000000011111111111100;
	memory[176] = 32'b00111111001111110011110000001111;
	memory[177] = 32'b00111100110011110011111111111111;
	memory[178] = 32'b00111100000011110011110000001111;
	memory[179] = 32'b00000000000000000011110000001111;
	memory[180] = 32'b00111111001111000011110000111100;
	memory[181] = 32'b00111111111111000011111111111100;
	memory[182] = 32'b00111100001111000011110011111100;
	memory[183] = 32'b00000000000000000011110000111100;
	memory[184] = 32'b00111100001111000000111111110000;
	memory[185] = 32'b00111100001111000011110000111100;
	memory[186] = 32'b00111100001111000011110000111100;
	memory[187] = 32'b00000000000000000000111111110000;
	memory[188] = 32'b00111100001111000011111111110000;
	memory[189] = 32'b00111111111100000011110000111100;
	memory[190] = 32'b00111100000000000011110000000000;
	memory[191] = 32'b00000000000000000011110000000000;
	memory[192] = 32'b00111100001111000000111111110000;
	memory[193] = 32'b00111100001111000011110000111100;
	memory[194] = 32'b00001111111100000011110000111100;
	memory[195] = 32'b00000000000000000000000011111100;
	memory[196] = 32'b00111100001111000011111111110000;
	memory[197] = 32'b00111111111100000011110000111100;
	memory[198] = 32'b00111100111100000011111111000000;
	memory[199] = 32'b00000000000000000011110000111100;
	memory[200] = 32'b00111100001111000000111111110000;
	memory[201] = 32'b00001111111100000011110000000000;
	memory[202] = 32'b00111100001111000000000000111100;
	memory[203] = 32'b00000000000000000000111111110000;
	memory[204] = 32'b00000011110000000011111111111100;
	memory[205] = 32'b00000011110000000000001111000000;
	memory[206] = 32'b00000011110000000000001111000000;
	memory[207] = 32'b00000000000000000000001111000000;
	memory[208] = 32'b00111100001111000011110000111100;
	memory[209] = 32'b00111100001111000011110000111100;
	memory[210] = 32'b00111100001111000011110000111100;
	memory[211] = 32'b00000000000000000000111111110000;
	memory[212] = 32'b00111100001111000011110000111100;
	memory[213] = 32'b00111100001111000011110000111100;
	memory[214] = 32'b00001111111100000011110000111100;
	memory[215] = 32'b00000000000000000000001111000000;
	memory[216] = 32'b00111100000011110011110000001111;
	memory[217] = 32'b00111100110011110011110000001111;
	memory[218] = 32'b00111111001111110011111111111111;
	memory[219] = 32'b00000000000000000011110000001111;
	memory[220] = 32'b00111100001111000011110000111100;
	memory[221] = 32'b00000011110000000000111111110000;
	memory[222] = 32'b00111100001111000000111111110000;
	memory[223] = 32'b00000000000000000011110000111100;
	memory[224] = 32'b00111100001111000011110000111100;
	memory[225] = 32'b00001111111100000011110000111100;
	memory[226] = 32'b00000011110000000000001111000000;
	memory[227] = 32'b00000000000000000000001111000000;
	memory[228] = 32'b00000000001111000011111111111100;
	memory[229] = 32'b00000011110000000000000011110000;
	memory[230] = 32'b00111100000000000000111100000000;
	memory[231] = 32'b00000000000000000011111111111100;
	memory[232] = 32'b00000000000000000000000000000000;
	memory[233] = 32'b00000000000000000000000000000000;
	memory[234] = 32'b00000011110000000000000000000000;
	memory[235] = 32'b00000000000000000000001111000000;
	memory[236] = 32'b00000000000000000000000000000000;
	memory[237] = 32'b00000000000000000000000000000000;
	memory[238] = 32'b00000011110000000000000000000000;
	memory[239] = 32'b00001111000000000000001111000000;
	memory[240] = 32'b00000000000000000000000000000000;
	memory[241] = 32'b00000000000000000000001111000000;
	memory[242] = 32'b00000011110000000000000000000000;
	memory[243] = 32'b00000000000000000000000000000000;
	memory[244] = 32'b00000000000000000000000000000000;
	memory[245] = 32'b00000000000000000000001111000000;
	memory[246] = 32'b00000011110000000000000000000000;
	memory[247] = 32'b00001111000000000000001111000000;
	memory[248] = 32'b00000000000000000000000000000000;
	memory[249] = 32'b00001111111111000000000000001111;
	memory[250] = 32'b00001111001111000011111100111100;
	memory[251] = 32'b00000000000000000000111100111100;
	memory[252] = 32'b00000011110000000000001111000000;
	memory[253] = 32'b00000011110000000000001111000000;
	memory[254] = 32'b00000000000000000000000000000000;
	memory[255] = 32'b00000000000000000000001111000000;
end

always@(posedge clk)
	out <= memory[addr[7:0]];

	
endmodule


